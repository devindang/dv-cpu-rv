//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2023, devin
//  balddonkey@outlook.com
//
//-------------------------------------------------------------------
// Title       : cpu_ctrl
// Author      : Devin
// Editor      : VIM
// Created     :
// Description :
//
// $Id$
//-------------------------------------------------------------------

`timescale 1ns / 1ps

module cpu_ctrl(
	input	
);


//------------------------ SIGNALS DECLARING GOES BELOW ------------------------//



//------------------------ PROCESS GOES BELOW ------------------------//



//------------------------ INSTANTIATE GOES BELOW ------------------------//


endmodule
