//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2023, devin
//  balddonkey@outlook.com
//
//-------------------------------------------------------------------
// Title       : rv_rf.V
// Author      : Devin
// Editor      : VIM
// Created     :
// Description :
//
// $Id$
//-------------------------------------------------------------------

`timescale 1ns / 1ps

module rv_rf(
    input   [4:0]   rd_reg1_i,
    input   [4:0]   rd_reg2_i,
    input   [4:0]   wr_reg_i,
    input   [63:0]  wr_data_i,
    output  [63:0]  rd_reg1_o,
    output  [63:0]  rd_reg2_o
);


//------------------------ SIGNALS ------------------------//



//------------------------ PROCESS ------------------------//



//------------------------ INST ------------------------//


endmodule