module rv_core(
    input clk,
);

endmodule