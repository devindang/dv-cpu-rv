module rv_data_path(
    input clk,
);

endmodule