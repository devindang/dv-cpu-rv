//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2023, devin
//  balddonkey@outlook.com
//
//-------------------------------------------------------------------
//
//  Author      : Devin
//  Project     : dv-cpu-rv
//  Repository  : https://github.com/devindang/dv-cpu-rv
//  Title       : rv_cpu_top.v
//  Dependances : rv_core
//  Editor      : code
//  Created     : 2023-08-24
//  Description : Process top design.
//
//-------------------------------------------------------------------

`timescale 1ns / 1ps

module rv_cpu_top(

);


//------------------------ SIGNALS ------------------------//



//------------------------ PROCESS ------------------------//



//------------------------ INST ------------------------//


endmodule